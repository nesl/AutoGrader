module MyWire(x, y);

	input wire x;
	output wire y;

	assign y = x;

endmodule

