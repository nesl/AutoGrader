module MyWire(dst_0, dst_1, src_1, src_0);
  output wire dst_0;
  output wire dst_1;
  input wire src_1;
  input wire src_0;
  assign dst_0 = src_0;
  assign dst_1 = src_1;
endmodule
